module instr_mem(input [31:0] addr, output [31:0] instr);
    reg [31:0] mem [0:255];
    initial $readmemh("instructions.mem", mem);
    assign instr = mem[addr];
endmodule